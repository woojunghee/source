library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
Library xpm;
use xpm.vcomponents.all;
use work.my_package.all;

entity ul_path_n77_100m is
port
(
    clk_491p52     : in  std_logic;
    clk_368p64     : in  std_logic;
    clk_122p88     : in  std_logic;
    clk_61p44      : in  std_logic;

    rst_n          : in  std_logic;

    tdd_sync       : in  std_logic;
    tsync_dly_in   : in std_logic_vector(1 downto 0);
    tsync_dly_out  : out arr_2_1_stdlogic;

    din_i          : in  arr_4_16_stdlogic;
    din_q          : in  arr_4_16_stdlogic;
    in_power       : out arr_4_32_stdlogic;
    in_peak        : out arr_4_32_stdlogic;
--    peak_sel       : in  std_logic;
--    pow_sel        : in  std_logic_vector(3 downto 0);

    input_gain     : in  arr_4_16_stdlogic;

    dc_path_en     : in  std_logic_vector(3 downto 0);
    dc_output_gain : in  arr_4_16_stdlogic;
    dc_out_pow     : out arr_4_32_stdlogic;
    dc_out_peak    : out arr_4_32_stdlogic;
    dc_dout_i      : out arr_4_16_stdlogic;
    dc_dout_q      : out arr_4_16_stdlogic;

    kd_path_en     : in  std_logic_vector(3 downto 0);
    kd_output_gain : in  arr_4_16_stdlogic;
    kd_out_pow     : out arr_4_32_stdlogic;
    kd_out_peak    : out arr_4_32_stdlogic;
    kd_dout_i      : out arr_4_16_stdlogic;
    kd_dout_q      : out arr_4_16_stdlogic;

    rm_path_en     : in  std_logic_vector(3 downto 0);
    rm_output_gain : in  arr_4_16_stdlogic;
    rm_out_pow     : out arr_4_32_stdlogic;
    rm_out_peak    : out arr_4_32_stdlogic;
    rm_dout_i      : out arr_4_16_stdlogic;
    rm_dout_q      : out arr_4_16_stdlogic;

    sb_path_en     : in  std_logic_vector(3 downto 0);
    sb_output_gain : in  arr_4_16_stdlogic;
    sb_out_pow     : out arr_4_32_stdlogic;
    sb_out_peak    : out arr_4_32_stdlogic;
    sb_dout_i      : out arr_4_16_stdlogic;
    sb_dout_q      : out arr_4_16_stdlogic;

    delay_dc_01    : in  std_logic_vector(13 downto 0);
    delay_dc_23    : in  std_logic_vector(13 downto 0);
    delay_kd_01    : in  std_logic_vector(13 downto 0);
    delay_kd_23    : in  std_logic_vector(13 downto 0);
    delay_rm_01    : in  std_logic_vector(13 downto 0);
    delay_rm_23    : in  std_logic_vector(13 downto 0);
    delay_sb_01    : in  std_logic_vector(13 downto 0);
    delay_sb_23    : in  std_logic_vector(13 downto 0);

    ul_iq_sync     : out std_logic

);
end ul_path_n77_100m;

architecture beh of ul_path_n77_100m is

----------------------------------------------------------------

  signal rst_n_122p88   : std_logic;
  signal rst_n_491p52   : std_logic;

  signal path_en        : std_logic_vector(MIMO_NUM downto 0);

  signal dc_dds         : std_logic_vector(31 downto 0);
  signal dc_dds_valid   : std_logic;
  signal kd_dds         : std_logic_vector(31 downto 0);
  signal kd_dds_valid   : std_logic;
  signal rm_dds         : std_logic_vector(31 downto 0);
  signal rm_dds_valid   : std_logic;
  signal sb_dds         : std_logic_vector(31 downto 0);
  signal sb_dds_valid   : std_logic;

  signal gain_out_i     : arr_mimo_16_stdlogic;
  signal gain_out_q     : arr_mimo_16_stdlogic;

  signal pow            : std_logic_vector(31 downto 0);

  signal dly_l_in       : std_logic_vector(31 downto 0);
  signal dly_l_out      : std_logic_vector(31 downto 0);

  signal fifo_empty     : std_logic;
  signal fifo_in        : std_logic_vector(31 downto 0);
  signal fifo_in_i      : std_logic_vector(15 downto 0);
  signal fifo_in_q      : std_logic_vector(15 downto 0);
  signal fifo_rd_en     : std_logic;
  signal fifo_in_valid  : std_logic;

  signal fifo_cnt       : integer range 0 to 1;

  signal cfr_in         : std_logic_vector(127 downto 0);
  signal cfr_in_valid   : std_logic;
  signal cfr_out        : std_logic_vector(127 downto 0);
  signal cfr_out_i      : arr_mimo_16_stdlogic;
  signal cfr_out_q      : arr_mimo_16_stdlogic;
  signal cfr_rdy        : std_logic;

  signal int2_in_i      : arr_mimo_16_stdlogic;
  signal int2_in_q      : arr_mimo_16_stdlogic;
  signal int2_in        : arr_mimo_32_stdlogic;
  signal int2_out_valid : std_logic_vector(MIMO_NUM downto 0);
  signal int2_out       : arr_mimo_128_stdlogic;


  signal dly_in_i       : std_logic_vector(15 downto 0);
  signal dly_in_q       : std_logic_vector(15 downto 0);
  signal dly_in         : std_logic_vector(31 downto 0);
  signal dly_out        : std_logic_vector(31 downto 0);
  signal dly_out_i      : std_logic_vector(15 downto 0);
  signal dly_out_q      : std_logic_vector(15 downto 0);

  signal dpd_in_buf_i   : std_logic_vector(15 downto 0);
  signal dpd_in_buf_q   : std_logic_vector(15 downto 0);

  signal gain_dout_i    : arr_mimo_16_stdlogic;
  signal gain_dout_q    : arr_mimo_16_stdlogic;

  signal pow_out_i      : std_logic_vector(15 downto 0);
  signal pow_out_q      : std_logic_vector(15 downto 0);
  signal pow_sel_s0     : std_logic_vector( 1 downto 0);
  signal pow_sel_s1     : std_logic_vector( 1 downto 0);
  signal out_pow        : std_logic_vector(31 downto 0);

  signal dc_off_ref     : std_logic_vector(15 downto 0) := x"0040";

  signal dc_det_i       : std_logic_vector(15 downto 0);
  signal dc_det_valid   : std_logic;

  signal dc_off_en      : std_logic;
  signal dc_off_en_s0   : std_logic;
  signal dc_off_en_s1   : std_logic;

  signal dc_off_in_i    : std_logic_vector(15 downto 0);
  signal dc_off_in_q    : std_logic_vector(15 downto 0);
  signal dc_off_out_i   : std_logic_vector(15 downto 0);
  signal dc_off_out_q   : std_logic_vector(15 downto 0);

  signal dc_din_i       : arr_4_16_stdlogic             := (others => (others => '0'));
  signal dc_din_q       : arr_4_16_stdlogic             := (others => (others => '0'));
  signal kd_din_i       : arr_4_16_stdlogic             := (others => (others => '0'));
  signal kd_din_q       : arr_4_16_stdlogic             := (others => (others => '0'));
  signal rm_din_i       : arr_4_16_stdlogic             := (others => (others => '0'));
  signal rm_din_q       : arr_4_16_stdlogic             := (others => (others => '0'));
  signal sb_din_i       : arr_4_16_stdlogic             := (others => (others => '0'));
  signal sb_din_q       : arr_4_16_stdlogic             := (others => (others => '0'));

  signal ul_iq_sync_cnt : std_logic_vector(1 downto 0);
  signal ul_iq_sync_s   : std_logic;
  signal rst_n_368p64   : std_logic;

  signal dc_user_in     : std_logic_vector(7 downto 0);
  signal dc_user_out    : std_logic_vector(7 downto 0);

  signal rm_user_in     : std_logic_vector(7 downto 0);
  signal rm_user_out    : std_logic_vector(7 downto 0);

attribute ASYNC_REG                   : string;
attribute ASYNC_REG of dc_off_en_s0   : signal is "true";
attribute ASYNC_REG of dc_off_en_s1   : signal is "true";


----------------------------------------------------------------
begin

rst_blk_122p88 : xpm_cdc_sync_rst
 generic map (
   DEST_SYNC_FF   => 2 ,
   INIT           => 1 ,
   INIT_SYNC_FF   => 0 ,
   SIM_ASSERT_CHK => 0 )
 port map (
   dest_rst       => rst_n_122p88 ,
   dest_clk       => clk_122p88   ,
   src_rst        => rst_n        );

rst_blk_368p64 : xpm_cdc_sync_rst
 generic map (
   DEST_SYNC_FF   => 2 ,
   INIT           => 1 ,
   INIT_SYNC_FF   => 0 ,
   SIM_ASSERT_CHK => 0 )
 port map (
   dest_rst       => rst_n_368p64 ,
   dest_clk       => clk_368p64   ,
   src_rst        => rst_n        );

rst_blk_491p52 : xpm_cdc_sync_rst
 generic map (
   DEST_SYNC_FF   => 2 ,
   INIT           => 1 ,
   INIT_SYNC_FF   => 0 ,
   SIM_ASSERT_CHK => 0 )
 port map (
   dest_rst       => rst_n_491p52 ,
   dest_clk       => clk_491p52   ,
   src_rst        => rst_n        );


in_pow_bank : for n in 0 to 3 generate
in_pow_mea : entity work.pow_mea_tdd_u
 generic map(
    clock_frequency => 491_520        , -- system clock frequency in khz 7_680, 15_360, 30_720, 61_440, 122_880, 245_760, 491_520
    unit_frequency  => 61_440         , -- unit clock frequency in khz 7_680, 5_760
    tdd_period      => 5_000          , -- tdd_period(us) 2_500, 5_000 ..
    tdd_high_time   => 1_142          , -- tdd_high_time(us) 3_857, 1_142
    check_time      => 20_000         ) -- check cycle(us) 20_000, 40_000, 80_000 ~ 320_000
 port map(
    clk             => clk_491p52     , --: in  std_logic;
    clk_unit        => clk_61p44      , --: in  std_logic;
    clk_tdd         => clk_122p88     , --: in  std_logic;
    reset_n         => rst_n_491p52   , --: in  std_logic;
    tdd_sync        => tdd_sync       , --: in  std_logic;
    din_i           => din_i(n)       , --: in  std_logic_vector(15 downto 0);
    din_q           => din_q(n)       , --: in  std_logic_vector(15 downto 0);
    din_vld         => '1'            , --: in  std_logic;
    chk_en          => '1'            , --: in  std_logic;
    power           => in_power(n)    , --: out std_logic_vector(31 downto 0);
    peak_power      => in_peak(n)     ); --: out std_logic_vector(31 downto 0)
end generate;

in_gain_bank : for n in 0 to mimo_num generate
in_gain_i : entity work.GAIN_BLK_16
 port map(
    clk     => clk_491p52     , --: in  std_logic;
    gain    => input_gain(n)  , --: in  std_logic_vector(15 downto 0);
    din     => din_i(n)       , --: in  std_logic_vector(15 downto 0);
    dout    => gain_out_i(n)  ); --: out std_logic_vector(15 downto 0)

in_gain_q : entity work.GAIN_BLK_16
 port map(
    clk     => clk_491p52     , --: in  std_logic;
    gain    => input_gain(n)  , --: in  std_logic_vector(15 downto 0);
    din     => din_q(n)       , --: in  std_logic_vector(15 downto 0);
    dout    => gain_out_q(n)  ); --: out std_logic_vector(15 downto 0)
end generate;


ul_dds_dcm : entity work.dds_dc_ul
port map
(
    aclk               => clk_491p52     , --: in std_logic;
    aresetn            => rst_n_491p52   , --: in std_logic;
    m_axis_data_tvalid => dc_dds_valid  , --: out std_logic;
    m_axis_data_tdata  => dc_dds        ); --: out std_logic_vector(31 downto 0);

ul_dds_kddi : entity work.dds_kd_ul
port map
(
    aclk               => clk_491p52     , --: in std_logic;
    aresetn            => rst_n_491p52   , --: in std_logic;
    m_axis_data_tvalid => kd_dds_valid , --: out std_logic;
    m_axis_data_tdata  => kd_dds       ); --: out std_logic_vector(31 downto 0);

ul_dds_rm : entity work.dds_rm_ul
port map
(
    aclk               => clk_491p52     , --: in std_logic;
    aresetn            => rst_n_491p52   , --: in std_logic;
    m_axis_data_tvalid => rm_dds_valid   , --: out std_logic;
    m_axis_data_tdata  => rm_dds         ); --: out std_logic_vector(31 downto 0);

ul_dds_sb : entity work.dds_sb_ul
port map
(
    aclk               => clk_491p52     , --: in std_logic;
    aresetn            => rst_n_491p52   , --: in std_logic;
    m_axis_data_tvalid => sb_dds_valid   , --: out std_logic;
    m_axis_data_tdata  => sb_dds         ); --: out std_logic_vector(31 downto 0);


ul_ddc_dc_bank : for n in 0 to mimo_num generate
ul_ddc_blk : entity work.ul_ddc
port map(
    clk_491p52          => clk_491p52        , --: in  std_logic;
    clk_122p88          => clk_122p88        , --: in  std_logic;
    clk_61p44           => clk_61p44         , --: in  std_logic;
    rst_n               => rst_n             , --: in  std_logic;
    din_i               => gain_out_i(n)     , --: in  std_logic_vector(15 downto 0);
    din_q               => gain_out_q(n)     , --: in  std_logic_vector(15 downto 0);
    tdd_sync            => tdd_sync          , --: in  std_logic;
    path_en             => dc_path_en(n)     , --: in  std_logic_vector(15 downto 0);
    dds_data            => dc_dds            , --: in  std_logic_vector(15 downto 0);
    dds_valid           => dc_dds_valid      , --: in  std_logic;
    output_gain         => dc_output_gain(n) , --: in  std_logic_vector(15 downto 0);
    out_pow             => dc_out_pow(n)     , --: out std_logic_vector(31 downto 0);
    out_peak            => dc_out_peak(n)    , --: out std_logic_vector(31 downto 0);
    dout_i              => dc_din_i(n)       , --: out std_logic_vector(15 downto 0);
    dout_q              => dc_din_q(n)       ); --: out std_logic_vector(15 downto 0)

end generate;

ul_ddc_kd_bank : for n in 0 to mimo_num generate
ul_ddc_blk : entity work.ul_ddc
port map(
    clk_491p52          => clk_491p52        , --: in  std_logic;
    clk_122p88          => clk_122p88        , --: in  std_logic;
    clk_61p44           => clk_61p44         , --: in  std_logic;
    rst_n               => rst_n             , --: in  std_logic;
    din_i               => gain_out_i(n)     , --: in  std_logic_vector(15 downto 0);
    din_q               => gain_out_q(n)     , --: in  std_logic_vector(15 downto 0);
    tdd_sync            => tdd_sync          , --: in  std_logic;
    path_en             => kd_path_en(n)     , --: in  std_logic_vector(15 downto 0);
    dds_data            => kd_dds            , --: in  std_logic_vector(15 downto 0);
    dds_valid           => kd_dds_valid      , --: in  std_logic;
    output_gain         => kd_output_gain(n) , --: in  std_logic_vector(15 downto 0);
    out_pow             => kd_out_pow(n)     , --: out std_logic_vector(31 downto 0);
    out_peak            => kd_out_peak(n)    , --: out std_logic_vector(31 downto 0);
    dout_i              => kd_din_i(n)       , --: out std_logic_vector(15 downto 0);
    dout_q              => kd_din_q(n)       ); --: out std_logic_vector(15 downto 0)

end generate;

ul_ddc_rm_bank : for n in 0 to mimo_num generate
ul_ddc_blk : entity work.ul_ddc
port map(
    clk_491p52          => clk_491p52        , --: in  std_logic;
    clk_122p88          => clk_122p88        , --: in  std_logic;
    clk_61p44           => clk_61p44         , --: in  std_logic;
    rst_n               => rst_n             , --: in  std_logic;
    din_i               => gain_out_i(n)     , --: in  std_logic_vector(15 downto 0);
    din_q               => gain_out_q(n)     , --: in  std_logic_vector(15 downto 0);
    tdd_sync            => tdd_sync          , --: in  std_logic;
    path_en             => rm_path_en(n)     , --: in  std_logic_vector(15 downto 0);
    dds_data            => rm_dds            , --: in  std_logic_vector(15 downto 0);
    dds_valid           => rm_dds_valid      , --: in  std_logic;
    output_gain         => rm_output_gain(n) , --: in  std_logic_vector(15 downto 0);
    out_pow             => rm_out_pow(n)     , --: out std_logic_vector(31 downto 0);
    out_peak            => rm_out_peak(n)    , --: out std_logic_vector(31 downto 0);
    dout_i              => rm_din_i(n)       , --: out std_logic_vector(15 downto 0);
    dout_q              => rm_din_q(n)         ); --: out std_logic_vector(15 downto 0)

end generate;

ul_ddc_sb_bank : for n in 0 to mimo_num generate
ul_ddc_blk : entity work.ul_ddc
port map(
    clk_491p52          => clk_491p52        , --: in  std_logic;
    clk_122p88          => clk_122p88        , --: in  std_logic;
    clk_61p44           => clk_61p44         , --: in  std_logic;
    rst_n               => rst_n             , --: in  std_logic;
    din_i               => gain_out_i(n)     , --: in  std_logic_vector(15 downto 0);
    din_q               => gain_out_q(n)     , --: in  std_logic_vector(15 downto 0);
    tdd_sync            => tdd_sync          , --: in  std_logic;
    path_en             => sb_path_en(n)     , --: in  std_logic_vector(15 downto 0);
    dds_data            => sb_dds            , --: in  std_logic_vector(15 downto 0);
    dds_valid           => sb_dds_valid      , --: in  std_logic;
    output_gain         => sb_output_gain(n) , --: in  std_logic_vector(15 downto 0);
    out_pow             => sb_out_pow(n)     , --: out std_logic_vector(31 downto 0);
    out_peak            => sb_out_peak(n)    , --: out std_logic_vector(31 downto 0);
    dout_i              => sb_din_i(n)       , --: out std_logic_vector(15 downto 0);
    dout_q              => sb_din_q(n)         ); --: out std_logic_vector(15 downto 0)

end generate;


dc_user_in(0)  <= tsync_dly_in(0);
tsync_dly_out(0)(0)   <= dc_user_out(0);

ul_dc_dly_blk0 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => dc_din_i(0)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => dc_din_q(0)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => dc_din_i(1)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => dc_din_q(1)  , --: in  std_logic_vector(15 downto 0);
    din_user        => dc_user_in   , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_dc_01  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => dc_dout_i(0) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => dc_dout_q(0) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => dc_dout_i(1) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => dc_dout_q(1) , --: out std_logic_vector(15 downto 0)
    dout_user       => dc_user_out  );--: out std_logic_vector(7 downto 0)

ul_dc_dly_blk1 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => dc_din_i(2)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => dc_din_q(2)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => dc_din_i(3)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => dc_din_q(3)  , --: in  std_logic_vector(15 downto 0);
    din_user        => x"00"        , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_dc_23  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => dc_dout_i(2) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => dc_dout_q(2) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => dc_dout_i(3) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => dc_dout_q(3) , --: out std_logic_vector(15 downto 0)
    dout_user       => open         );--: out std_logic_vector(7 downto 0)


ul_kd_dly_blk0 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => kd_din_i(0)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => kd_din_q(0)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => kd_din_i(1)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => kd_din_q(1)  , --: in  std_logic_vector(15 downto 0);
    din_user        => x"00"        , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_kd_01  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => kd_dout_i(0) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => kd_dout_q(0) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => kd_dout_i(1) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => kd_dout_q(1) , --: out std_logic_vector(15 downto 0)
    dout_user       => open         );--: out std_logic_vector(7 downto 0)

ul_kd_dly_blk1 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => kd_din_i(2)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => kd_din_q(2)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => kd_din_i(3)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => kd_din_q(3)  , --: in  std_logic_vector(15 downto 0);
    din_user        => x"00"        , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_kd_23  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => kd_dout_i(2) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => kd_dout_q(2) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => kd_dout_i(3) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => kd_dout_q(3) , --: out std_logic_vector(15 downto 0)
    dout_user       => open         );--: out std_logic_vector(7 downto 0)

rm_user_in(0)    <= tsync_dly_in(1);
tsync_dly_out(1)(0) <= rm_user_out(0);

ul_rm_dly_blk0 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => rm_din_i(0)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => rm_din_q(0)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => rm_din_i(1)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => rm_din_q(1)  , --: in  std_logic_vector(15 downto 0);
    din_user        => rm_user_in   , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_rm_01  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => rm_dout_i(0) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => rm_dout_q(0) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => rm_dout_i(1) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => rm_dout_q(1) , --: out std_logic_vector(15 downto 0)
    dout_user       => rm_user_out  );--: out std_logic_vector(7 downto 0)

ul_rm_dly_blk1 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => rm_din_i(2)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => rm_din_q(2)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => rm_din_i(3)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => rm_din_q(3)  , --: in  std_logic_vector(15 downto 0);
    din_user        => x"00"        , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_rm_23  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => rm_dout_i(2) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => rm_dout_q(2) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => rm_dout_i(3) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => rm_dout_q(3) , --: out std_logic_vector(15 downto 0)
    dout_user       => open         );--: out std_logic_vector(7 downto 0)

ul_sb_dly_blk0 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => sb_din_i(0)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => sb_din_q(0)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => sb_din_i(1)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => sb_din_q(1)  , --: in  std_logic_vector(15 downto 0);
    din_user        => x"00"        , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_sb_01  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => sb_dout_i(0) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => sb_dout_q(0) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => sb_dout_i(1) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => sb_dout_q(1) , --: out std_logic_vector(15 downto 0)
    dout_user       => open         );--: out std_logic_vector(7 downto 0)

ul_sb_dly_blk1 : entity work.delay_blk_uram
port map(
    clk             => clk_122p88   , --: in  std_logic;
    rst_n           => rst_n        , --: in  std_logic;
    din_i_m0        => sb_din_i(2)  , --: in  std_logic_vector(15 downto 0);
    din_q_m0        => sb_din_q(2)  , --: in  std_logic_vector(15 downto 0);
    din_i_m1        => sb_din_i(3)  , --: in  std_logic_vector(15 downto 0);
    din_q_m1        => sb_din_q(3)  , --: in  std_logic_vector(15 downto 0);
    din_user        => x"00"        , --: in  std_logic_vector(7 downto 0);
    delay_parameter => delay_sb_23  , --: in  std_logic_vector(13 downto 0);
    dout_i_m0       => sb_dout_i(2) , --: out std_logic_vector(15 downto 0);
    dout_q_m0       => sb_dout_q(2) , --: out std_logic_vector(15 downto 0);
    dout_i_m1       => sb_dout_i(3) , --: out std_logic_vector(15 downto 0);
    dout_q_m1       => sb_dout_q(3) , --: out std_logic_vector(15 downto 0)
    dout_user       => open         );--: out std_logic_vector(7 downto 0)

process(clk_368p64)
begin
if rising_edge(clk_368p64) then
    if (rst_n_368p64 = '0') then
        ul_iq_sync_cnt <= "00";
    else
        if (ul_iq_sync_cnt = "10") then
            ul_iq_sync_cnt <= "00";
        else
            ul_iq_sync_cnt <= ul_iq_sync_cnt+1;
        end if;
    end if;
end if;
end process;

process(clk_368p64)
begin
if rising_edge(clk_368p64) then
    if (ul_iq_sync_cnt = "01") then
        ul_iq_sync_s <= '1';
    else
        ul_iq_sync_s <= '0';
    end if;
end if;
end process;

ul_iq_sync <= ul_iq_sync_s;


end beh;

